library verilog;
use verilog.vl_types.all;
entity seven_seg_B_tm is
end seven_seg_B_tm;
