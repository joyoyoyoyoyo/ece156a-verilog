module dff_B(clk, q, q_bar, d);
  output q, q_bar;
  input clk, d;
  
  always @ (posedge clk)
  begin
      
  end
endmodule
    
