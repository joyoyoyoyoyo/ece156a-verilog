library verilog;
use verilog.vl_types.all;
entity dff_B_tm is
end dff_B_tm;
